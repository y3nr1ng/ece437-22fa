`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/25/2022 01:28:42 PM
// Design Name: 
// Module Name: drv8833
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module drv8833 #(
    parameter PULSE_CLK_DIVIDER = 16'd250 
)(
    input               i_clk, 
    
    // control
    input               i_rst,
    input               i_start,
    
    input               i_dir,
    input       [23:0]  i_pulses,
    
    output reg          o_done,
    
    // wirings
    output              o_pmod_dir,
    output              o_pmod_en
);
    
    /*** en pulse generator ***/
    reg [15:0]  pmod_en_counter = 0;
    reg         pmod_en = 0;
    
    always @(posedge i_clk) begin
        if (i_rst) begin
            pmod_en_counter <= 0;
        end
        else begin
            if (pmod_en_counter >= PULSE_CLK_DIVIDER/2) begin
                pmod_en_counter <= 0;
                pmod_en <= ~pmod_en;
            end
            else begin
                pmod_en_counter <= pmod_en_counter + 1'b1;
            end
        end
    end
    
    reg pmod_oe = 0; // this is what we want to control 
    assign o_pmod_en = (pmod_oe & !i_rst) & pmod_en;
    
    wire pmod_en_tick;
    assign pmod_en_tick = (pmod_en_counter == PULSE_CLK_DIVIDER/2) & o_pmod_en;
    /*** en pulse generator ***/
    
    /*** en counter ***/
    reg         clear = 0;
    reg [23:0]  counter = 0;
    
    always @(posedge pmod_en or posedge clear) begin
        if (clear) begin
            counter <= 0;
        end
        else begin
            counter <= counter + 1'b1;
        end
    end
    /*** en counter ***/
    
    /*** dir control ***/
    reg dir = 0;
    assign o_pmod_dir = dir;
    /*** dir control ***/
    
    /*** main fsm ***/
    integer state;
    localparam S_IDLE = 0,
               S_PREPARE = 1,
               S_RUN = 2;
    
    reg start = 0;

    reg [23:0] target_counter = 0;
    
    always @(posedge i_clk) begin
        o_done <= 0;
        if (o_done) begin
            start <= 0;
        end

        if (i_start) begin
            start <= 1;
        end
        
        if (i_rst) begin 
            state <= S_IDLE;
         
            // dir and en
            dir <= 0;
            pmod_oe <= 0;
            
            // en counter
            clear <= 1;
            target_counter <= 0;   
        end 
        else begin
            

            case (state)
                S_IDLE: begin
                    if (start) begin
                        state <= S_PREPARE;
                    end
                end

                S_PREPARE: begin
                    // set_direction
                    dir <= i_dir;

                    // reset pulse counter 
                    clear <= 1;
                    target_counter <= i_pulses;

                    pmod_oe <= 1;

                    state <= S_RUN;
                end
                
                S_RUN: begin
                    clear <= 0;
                    
                    if (counter >= target_counter) begin
                        pmod_oe <= 0;
                        o_done <= 1;
                        state <= S_IDLE;
                    end
                end
            endcase
        end
    end
    
    assign o_busy = (state != S_IDLE);
    /*** main fsm ***/
    
endmodule
